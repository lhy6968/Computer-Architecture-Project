`timescale 1ns/1ps

// general register
`define gr0  	5'b00000
`define gr1  	5'b00001
`define gr2  	5'b00010
`define gr3 	5'b00011
`define gr4  	5'b00100
`define gr5  	5'b00101
`define gr6  	5'b00110
`define gr7  	5'b00111
`define gr8  	5'b01000
`define gr9  	5'b01001
`define gr10  	5'b01010
`define gr11  	5'b01011
`define gr12  	5'b01100
`define gr13  	5'b01101
`define gr14  	5'b01110
`define gr15  	5'b01111
`define gr16  	5'b10000
`define gr17  	5'b10001
`define gr18  	5'b10010
`define gr19  	5'b10011
`define gr20  	5'b10100
`define gr21  	5'b10101
`define gr22  	5'b10110
`define gr23 	5'b10111
`define gr24  	5'b11000
`define gr25  	5'b11001
`define gr26  	5'b11010
`define gr27  	5'b11011
`define gr28  	5'b11100
`define gr29  	5'b11101
`define gr30  	5'b11110
`define gr31  	5'b11111

module CPU_test;

    // Inputs
	reg clock;
	reg [31:0] d_datain;
	reg [31:0] i_datain;
    reg start;

    wire [31:0] d_dataout;
    wire [31:0] d_addr;

    CPU uut(
        .clock(clock),
        .start(start), 
		.d_datain(d_datain), 
		.i_datain(i_datain),
        .d_dataout(d_dataout),
        .d_addr(d_addr)
    );

    initial begin
        // Initialize Inputs
        clock = 0;
        start = 1;

    $display("pc  :        instruction             :  gr0   :  gr1   :  gr2   :  gr3   :   gr31 :dataout : address");
    $monitor("%h:%b:%h:%h:%h:%h:%h:%h:%h", 
        uut.pc,i_datain, uut.gr[0], uut.gr[1], uut.gr[2], uut.gr[3],uut.gr[31],d_dataout,d_addr);

    /*Test:*/
//lw
    #period
    d_datain <= 32'h0000_00ab;
    i_datain <= {6'b100011, `gr0, `gr1, 16'h0001};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//lw
    #period d_datain <= 32'h0000_3c00;
    i_datain <= {6'b100011, `gr0, `gr2, 16'h0002};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;


//add
    #period i_datain <= {6'b000000, `gr1, `gr2, `gr3,  5'b00000, 6'b100000};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;


//addu
    #period i_datain <= {6'b000000, `gr2, `gr3, `gr1,  5'b00000, 6'b100001};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//addi
    #period i_datain <= {6'b001000,`gr3, `gr1,  16'b0000000000001000};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//addiu
    #period i_datain <= {6'b001001,`gr2, `gr1,  16'b0000000000001001};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//sub
    #period i_datain <= {6'b000000, `gr1, `gr2, `gr3,  5'b00000, 6'b100010};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//subu
    #period i_datain <= {6'b000000, `gr2, `gr3, `gr1,  5'b00000, 6'b100011};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//and
    #period i_datain <= {6'b000000, `gr1, `gr2, `gr3,  5'b00000, 6'b100100};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//andi
    #period i_datain <= {6'b001100,`gr2, `gr1,  16'b1110000000001111};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//or
    #period i_datain <= {6'b000000, `gr1, `gr2, `gr3,  5'b00000, 6'b100101};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//ori
    #period i_datain <= {6'b001101,`gr2, `gr1,  16'b1110000000011111};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//nor
    #period i_datain <= {6'b000000, `gr1, `gr2, `gr3,  5'b00000, 6'b100111};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//xor
    #period i_datain <= {6'b000000, `gr1, `gr2, `gr3,  5'b00000, 6'b100110};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//sll
    #period i_datain <= {6'b000000, `gr1, `gr2, `gr3,  5'b00010, 6'b000000};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//sra
    #period i_datain <= {6'b000000, `gr1, `gr2, `gr3,  5'b00010, 6'b000011};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//srl
    #period i_datain <= {6'b000000, `gr2, `gr1, `gr3,  5'b00011, 6'b000010};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//lw
    #period d_datain <= 32'b00000000000000000000000000000011;
    i_datain <= {6'b100011, `gr0, `gr2, 16'h0002};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//sllv
    #period i_datain <= {6'b000000, `gr2, `gr3, `gr1,  5'b00000, 6'b000100};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//srav
    #period i_datain <= {6'b000000, `gr2, `gr1, `gr3,  5'b00000, 6'b000111};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//srlv
    #period i_datain <= {6'b000000, `gr2, `gr3, `gr1,  5'b00000, 6'b000110};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//slt
    #period i_datain <= {6'b000000, `gr3, `gr2, `gr1,  5'b00000, 6'b101010};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//jr
    #period i_datain <= {6'b000000, `gr2,21'b000000000000000001000};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//j
    #period i_datain <= {6'b000010, 26'b00000000000011111111111111};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//jal
    #period i_datain <= {6'b000011, 26'b00000000000011111111110000};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//beq
    #period i_datain <= {6'b000100,`gr0,`gr0,16'b0000000000001111};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
//bne
    #period i_datain <= {6'b000101,`gr0,`gr0,16'b0000000000001111};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;


    #period i_datain <= {6'b000000, `gr3, `gr2, `gr1,  5'b00000, 6'b100000};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

//sw
    #period i_datain <= {6'b101011,`gr0,`gr1,16'b0000000000001111};
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    #period i_datain <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;




    #period $finish;
    end

parameter period = 10;
always #5 clock = ~clock;
endmodule