`timescale 1ns/1ps

module alu_test;

reg[31:0] i_datain,gr1,gr2;

wire[31:0]hi;
wire[31:0]lo;
wire[31:0]c;
wire[2:0]zon;


alu testalu(i_datain,gr1,gr2,c,zon,hi,lo);

initial
begin


$display("instruction:op:func:  gr1   :   gr2  : reg_A  : reg_B  : reg_C  :   lo   :   hi   :zon");
$monitor("   %h:%h: %h :%h:%h:%h:%h:%h:%h:%h:%b",
i_datain, testalu.opcode, testalu.func, gr1 , gr2, testalu.reg_A, testalu.reg_B, testalu.reg_C,testalu.reg_lo,testalu.reg_hi,zon);

//// arith left shift
//add
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
gr2 <=32'b1101_1101_1101_1101_1101_1101_1101_1101;
//addi
#10 i_datain<=32'b0010_0000_0000_0000_1111_1111_1111_1111;
gr1 <=32'b0111_1111_1111_1111_1111_1111_1111_1111;
//addu
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
gr1 <=32'b0100_0000_0100_0000_0100_0000_0100_0000;
gr2 <=32'b0101_1101_1101_1101_1101_1101_1101_1101;
//addiu
#10 i_datain<=32'b0010_0100_0000_0001_1111_1111_1111_1111;
gr1 <=32'b0100_0000_0100_0000_0100_0000_0100_0000;
//sub
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
gr1 <=32'b0101_1101_1101_1101_1101_1101_1101_1101;
gr2 <=32'b0101_1101_1101_1101_1101_1101_1101_1101;
//subu
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
gr1 <=32'b0111_1111_1111_1111_1111_1111_1111_1111;
gr2 <=32'b0000_0000_0000_0000_1111_1111_1111_1111;
//mult
#10 i_datain<=32'b0000_0000_0000_0001_0000_0000_0001_1000;
gr1 <=32'b1111_1111_1111_1111_1111_1111_1111_1111;
gr2 <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
//multu
#10 i_datain<=32'b0000_0000_0000_0001_0000_0000_0001_1001;
gr1 <=32'b0000_0000_0000_0000_0000_0000_0000_1101;
gr2 <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
//div
#10 i_datain<=32'b0000_0000_0000_0001_0000_0000_0001_1010;
gr1 <=32'b1111_1111_1111_1111_1111_1111_1110_0001;
gr2 <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
//divu
#10 i_datain<=32'b0000_0000_0000_0001_0000_0000_0001_1011;
gr1 <=32'b0000_0000_0000_0000_0000_0000_0000_1101;
gr2 <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
//and
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0100;
gr1<=32'b1111_1111_1111_1111_1111_1111_1111_0001;
gr2 <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
//andi
#10 i_datain<=32'b0011_0000_0100_0001_0000_0000_0001_0001;
gr1<=32'b1111_1111_1111_1111_1111_1111_1110_0001;
//or
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0101;
gr1<=32'b0101_1001_1101_1101_1101_0001_1101_1101;
gr2 <=32'b0111_1001_1101_1101_1101_0001_1101_1101;
//ori
#10 i_datain<=32'b0011_0100_0100_0001_0000_0000_0001_0001;
gr1<=32'b1111_1111_1111_1111_1111_1111_1110_0001;
//nor
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0111;
gr1<=32'b1111_1111_1111_1111_1111_1111_1110_0001;
gr2 <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
//xor
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0110;
gr1<=32'b1111_1111_1111_1111_1111_1111_1110_0001;
gr2 <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
//xori
#10 i_datain<=32'b0011_1000_0100_0001_0000_0000_0001_0001;
gr1<=32'b1111_1111_1111_1111_1111_1111_1110_0001;
//beq
#10 i_datain<=32'b0001_0000_0000_0001_0000_0000_0010_0000;
gr1 <=32'b0101_1101_1101_1101_1101_1101_1101_1101;
gr2 <=32'b0101_1101_1101_1101_1101_1101_1101_1101;
//slt
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
gr2 <=32'b1101_1101_1101_1101_1101_1101_1101_1101;
//slti
#10 i_datain<=32'b0010_1000_0100_0001_0000_0000_0000_1101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
//bne
#10 i_datain<=32'b0001_0100_0000_0001_0000_0000_0010_0000;
gr1 <=32'b0101_1101_1101_1101_1101_1101_1101_1101;
gr2 <=32'b0101_1101_1101_1101_1101_1101_1101_1101;
//sltu
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
gr2 <=32'b1101_1101_1101_1101_1101_1101_1101_1101;
//sltiu
#10 i_datain<=32'b0010_1100_0100_0001_0000_0000_0000_1101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
//lw
#10 i_datain<=32'b1000_1100_0100_0001_0000_0000_0010_0000;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
gr2 <=32'b1101_1101_1101_1101_1101_1101_1101_1101;
//sll
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0000;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
//sllv
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0100;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
//srl
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0010;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
//srlv
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0110;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
//sw
#10 i_datain<=32'b1010_1110_0000_0001_0000_0000_0010_0000;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
gr2 <=32'b1101_1101_1101_1101_1101_1101_1101_1101;
//sra
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0011;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
//srav
#10 i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0111;
gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;


#10 $finish;
end

endmodule