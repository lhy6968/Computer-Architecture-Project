
`timescale 1ns/1ps
module alu_test;

reg[31:0] a,b;
reg[5:0] opcode;

wire[31:0] hi;
wire[31:0] lo;
wire[31:0] c;
wire zero;
wire overflow;
wire neg;
wire[2:0] zon;


parameter  add = 6'b000001,
addi = 6'b000010,
addu = 6'b000011,
addiu = 6'b000100,
sub  = 6'b000101,
subu  = 6'b000110,
mult = 6'b000111,
multu  = 6'b001000,
div = 6'b001001,
divu = 6'b001010,
sqrt = 6'b001011,
and_ = 6'b001100,
andi = 6'b001101,
or_ = 6'b001110,
ori  = 6'b001111,
nor_ = 6'b010000,
xor_  = 6'b010001,
xnor_ = 6'b010010, 
slt = 6'b010011,
slti = 6'b010100;


alu testalu(a,b,opcode,c,zon,hi,lo);


initial
begin

$display("op: a      : b      : c      : hi      :lo      :   zon");
$monitor(" %h:%h:%h:%h:%h:%h:%b",
opcode, a, b, c, hi, lo, zon);

//// arith left shift



#10 a=32'b0100_0000_0100_0000_0100_0000_0100_0000;
b = 32'b1101_1101_1101_1101_1101_1101_1101_1101;
opcode= add;

#10 a=32'b0100_0000_0100_0000_0100_0000_0100_0000;
b = 32'b0101_1101_1101_1101_1101_1101_1101_1101;
opcode= add;

#10 a=32'b0111_1111_1111_1111_1111_1111_1111_1111;
b = 32'b0000_0000_0000_0000_1111_1111_1111_1111;
opcode= addi;

#10 a=32'b0100_0000_0100_0000_0100_0000_0100_0000;
b = 32'b0101_1101_1101_1101_1101_1101_1101_1101;
opcode= addu;

#10 a=32'b0100_0000_0100_0000_0100_0000_0100_0000;
b = 32'b0000_0000_0000_0000_1111_1111_1111_1111;
opcode= addiu;

#10 a=32'b0101_1101_1101_1101_1101_1101_1101_1101;
b = 32'b0101_1101_1101_1101_1101_1101_1101_1101;
opcode= sub;

#10 a=32'b0111_1111_1111_1111_1111_1111_1111_1111;
b = 32'b0000_0000_0000_0000_1111_1111_1111_1111;
opcode= subu;

#10 a=32'b1111_1111_1111_1111_1111_1111_1111_1111;
b = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
opcode= mult;
#10 a=32'b0000_0000_0000_0000_0000_0000_0000_1101;
b = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
opcode= multu;


#10 a=32'b1111_1111_1111_1111_1111_1111_1110_0001;
b = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
opcode= div;

#10 a=32'b0000_0000_0000_0000_0000_0000_0000_1101;
b = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
opcode= divu;

#10 a=32'b0000_0000_0000_0000_0000_0000_0111_1010;
b = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
opcode= sqrt;

#10 a=32'b1111_1111_1111_1111_1111_1111_1111_0001;
b = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
opcode = and_ ;

#10 a=32'b1111_1111_1111_1111_1111_1111_1110_0001;
b = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
opcode= andi;

#10 a=32'b0101_1001_1101_1101_1101_0001_1101_1101;
b = 32'b0111_1001_1101_1101_1101_0001_1101_1101;
opcode= or_;

#10 a=32'b1111_1111_1111_1111_1111_1111_1110_0001;
b = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
opcode= ori;

#10 a=32'b1111_1111_1111_1111_1111_1111_1110_0001;
b = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
opcode= nor_;

#10 a=32'b1111_1111_1111_1111_1111_1111_1110_0001;
b = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
opcode= xor_;

#10 a=32'b1111_1111_1111_1111_1111_1111_1110_0001;
b = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
opcode= xnor_;


#10 a=32'b1101_1101_1101_1101_1101_1101_1101_1100;
b = 32'b1101_1101_1101_1101_1101_1101_1101_1101;
opcode= slt;

#10 a=32'b0100_0000_0100_0000_0100_0000_0100_0000;
b = 32'b1101_1101_1101_1101_1101_1101_1101_1101;
opcode= slt;
#10 a=32'b0000_0000_0000_0000_0000_0000_0000_0001;
b = 32'b0000_0000_0000_0000_0000_0000_0000_1101;
opcode= slti;
#10 $finish;
end
endmodule


